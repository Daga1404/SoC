`timescale 1ns/1ps

module main_decoder_tb;
    // Inputs
    reg clk;
    reg [6:0] op;
    
    // Outputs
    wire branch;
    wire jump;
    wire mem_write;
    wire alu_src;
    wire reg_write;
    wire [1:0] result_src;
    wire [1:0] imm_src;
    wire [1:0] alu_op;
    
    // Instantiate the Unit Under Test (UUT)
    main_decoder uut (
        .clk(clk),
        .op(op),
        .branch(branch),
        .jump(jump),
        .mem_write(mem_write),
        .alu_src(alu_src),
        .reg_write(reg_write),
        .result_src(result_src),
        .imm_src(imm_src),
        .alu_op(alu_op)
    );
    
    // Clock generation
    always #5 clk = ~clk;
    
    // Test case checker
    task check_outputs;
        input expected_branch;
        input expected_jump;
        input expected_mem_write;
        input expected_alu_src;
        input expected_reg_write;
        input [1:0] expected_result_src;
        input [1:0] expected_imm_src;
        input [1:0] expected_alu_op;
        input [6:0] opcode;
        begin
            if (branch !== expected_branch) $display("ERROR at opcode %d: branch = %b, expected %b", opcode, branch, expected_branch);
            if (jump !== expected_jump) $display("ERROR at opcode %d: jump = %b, expected %b", opcode, jump, expected_jump);
            if (mem_write !== expected_mem_write) $display("ERROR at opcode %d: mem_write = %b, expected %b", opcode, mem_write, expected_mem_write);
            if (alu_src !== expected_alu_src && expected_alu_src !== 1'bx) $display("ERROR at opcode %d: alu_src = %b, expected %b", opcode, alu_src, expected_alu_src);
            if (reg_write !== expected_reg_write) $display("ERROR at opcode %d: reg_write = %b, expected %b", opcode, reg_write, expected_reg_write);
            if (result_src !== expected_result_src && expected_result_src !== 2'bxx) $display("ERROR at opcode %d: result_src = %b, expected %b", opcode, result_src, expected_result_src);
            if (imm_src !== expected_imm_src && expected_imm_src !== 2'bxx) $display("ERROR at opcode %d: imm_src = %b, expected %b", opcode, imm_src, expected_imm_src);
            if (alu_op !== expected_alu_op && expected_alu_op !== 2'bxx) $display("ERROR at opcode %d: alu_op = %b, expected %b", opcode, alu_op, expected_alu_op);
            $display("Test case for opcode %d completed", opcode);
        end
    endtask
    
    initial begin
        // Initialize inputs
        clk = 0;
        op = 0;
        
        // Wait for global reset
        #20;
        
        // Test case 1: Load Word (lw) - op = 3
        op = 7'd3;
        #15; // Wait for clock edge and some settling time
        check_outputs(
            1'b0,    // branch
            1'b0,    // jump
            1'b0,    // mem_write
            1'b1,    // alu_src
            1'b1,    // reg_write
            2'b01,   // result_src
            2'b00,   // imm_src
            2'b00,   // alu_op
            7'd3     // opcode for reference
        );
        
        // Test case 2: I-Type - op = 19
        op = 7'd19;
        #10; // One clock cycle
        check_outputs(
            1'b0,    // branch
            1'b0,    // jump
            1'b0,    // mem_write
            1'b1,    // alu_src
            1'b1,    // reg_write
            2'b00,   // result_src
            2'b00,   // imm_src
            2'b10,   // alu_op
            7'd19    // opcode for reference
        );
        
        // Test case 3: R-Type - op = 51
        op = 7'd51;
        #10;
        check_outputs(
            1'b0,    // branch
            1'b0,    // jump
            1'b0,    // mem_write
            1'b0,    // alu_src
            1'b1,    // reg_write
            2'b00,   // result_src
            2'bxx,   // imm_src (don't care)
            2'b10,   // alu_op
            7'd51    // opcode for reference
        );
        
        // Test case 4: Store Word (sw) - op = 35
        op = 7'd35;
        #10;
        check_outputs(
            1'b0,    // branch
            1'b0,    // jump
            1'b1,    // mem_write
            1'b1,    // alu_src
            1'b0,    // reg_write
            2'bxx,   // result_src (don't care)
            2'b01,   // imm_src
            2'b00,   // alu_op
            7'd35    // opcode for reference
        );
        
        // Test case 5: Branch Equal (beq) - op = 99
        op = 7'd99;
        #10;
        check_outputs(
            1'b1,    // branch
            1'b0,    // jump
            1'b0,    // mem_write
            1'b0,    // alu_src
            1'b0,    // reg_write
            2'bxx,   // result_src (don't care)
            2'b01,   // imm_src
            2'b01,   // alu_op
            7'd99    // opcode for reference
        );
        
        // Test case 6: Jump and Link (jal) - op = 111
        op = 7'd111;
        #10;
        check_outputs(
            1'b0,    // branch
            1'b1,    // jump
            1'b0,    // mem_write
            1'bx,    // alu_src (don't care)
            1'b1,    // reg_write
            2'b10,   // result_src
            2'b11,   // imm_src
            2'bxx,   // alu_op (don't care)
            7'd111   // opcode for reference
        );
        
        // Test case 7: Default case - op = 0
        op = 7'd0;
        #10;
        check_outputs(
            1'b0,    // branch
            1'b0,    // jump
            1'b0,    // mem_write
            1'b0,    // alu_src
            1'b0,    // reg_write
            2'b00,   // result_src
            2'b00,   // imm_src
            2'b00,   // alu_op
            7'd0     // opcode for reference
        );
        
        // Test case 8: Another invalid opcode
        op = 7'd127;
        #10;
        check_outputs(
            1'b0,    // branch
            1'b0,    // jump
            1'b0,    // mem_write
            1'b0,    // alu_src
            1'b0,    // reg_write
            2'b00,   // result_src
            2'b00,   // imm_src
            2'b00,   // alu_op
            7'd127   // opcode for reference
        );
        
        $display("All tests completed");
        //#10 $finish;
    end
    
    // Optional: Dump waveform to a VCD file for viewing in a waveform viewer
    initial begin
        $dumpfile("main_decoder_tb.vcd");
        $dumpvars(0, main_decoder_tb);
    end
    
endmodule